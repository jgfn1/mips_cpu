module Shift_left2(input[31:0] S_end, output[31:0] saida32);


		always_comb
			begin 
				saida32 =(S_ent << 2)			
			
			end
		
		endmodule
		
		
		