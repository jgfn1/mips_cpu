module mux32_2_1 (input logic )